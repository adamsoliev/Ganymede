/* verilator lint_off UNUSED */
module CPU(input    logic   clk_i);
        
    // logic [12:0] counter;
    // always @(posedge clk_i) begin
    //     counter <= counter + 1;
    // end

    // assign led_o = counter[11];

endmodule
/* verilator lint_off UNUSED */